module usr(
		input clk,
		input [1:0]sel,
		input [3:0]ip,
		input leftS,
		input rightS,

		output [3:0]q,
		output [3:0]qb,
		output [3:0]y	);


demux dm0	( sel, {ip[3], q[2], rightS, q[3]}, y[3]   );
d_ff d0		( y[3], clk, q[3], qb[3] );

demux dm1	( sel, {ip[2], q[1], q[3], q[2]}, y[2]   );
d_ff d1		( y[2], clk, q[2], qb[2] );

demux dm2	( sel, {ip[1], q[0], q[2], q[1]}, y[1]   );
d_ff d2		( y[1], clk, q[1], qb[1] );

demux dm3	( sel, {ip[0], leftS, q[1], q[0]}, y[1]   );
d_ff d3		( y[0], clk, q[0], qb[0] );


endmodule


module demux(
		input [1:0]sel,
		input [3:0]ip,

		output reg y	);

always @(sel)
begin
	case(sel)
	
	2'b00:  y	=	ip[0];	// No changes
	2'b01:	y	=	ip[1];	// Right Shift
	2'b10:	y	=	ip[2];	// Left Shift 
	2'b11:	y	=	ip[3];	// Parallel Input 

	endcase
end

endmodule


module d_ff(
		input d,
		input clk,
		
		output reg q,
		output reg qb	);

always @(posedge clk)
begin
	q 	=	 d;	
	qb	=	~q;
end

endmodule

