module bin2xs3(

		input [3:0]bin,
		output [3:0]xs3
				);

assign xs3 = bin + 4'd3;

// assign xs3 = bin + 4'b0011;

endmodule


