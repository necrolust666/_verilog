
/* 
Design
*/

module halfAdder(val1, val2, sum, carry);
  
  	input wire val1, val2;
  	output reg sum, carry;
  
/*
 	// Gate Level/Structural Modelling
  
	xor(sum, val1, val2);
	and(carry, val1, val2);
*/
 
/*
	// Data Flow Modelling/RTL Level Modelling/Conditional Modelling
	assign sum = val1^val2;
	assign carry = val1&val2;
*/

	// Behavorial Modelling	
	always @(*)	// * == Any Event
	begin
/*		
	case({val1, val2})

	2'b00: begin sum=1'b0; carry=1'b0; end
	2'b01: begin sum=1'b1; carry=1'b0; end
	2'b10: begin sum=1'b1; carry=1'b0; end
	2'b11: begin sum=1'b0; carry=1'b1; end
	endcase
*/
	assign {carry, sum} = val1 + val2;
	end

endmodule
